`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/03/2023 09:33:38 PM
// Design Name: 
// Module Name: crc7
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module crc7
(
    input clk_i,
    input rst_i,
    input en_i,
    input [39:0] data_i
    output [6:0] crc_o,
    output crc_valid_o
);


endmodule
